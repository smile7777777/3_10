** 111062307_HW1 **
** Environment setting **
*************************
*      Your code        *
*************************

*** Inverter ***
.subckt INV in1 inv_out vdd vss
** Your code **
.ends

*** OR ***
.subckt OR2 in2 in3 OR vdd vss
** Your code **
.ends

*** AND ***
.subckt AND2 in4 in5 AND vdd vss
** Your code **
.ends

*** logic function ***
.subckt logic A B C D F vdd vss
** Your code **
.ends