** 123456_HW1_bonus **
** Environment setting **
*************************
*      Your code        *
*************************

*** 4 to 1 MUX ***
.subckt MUX S0 S1 D0 D1 D2 D3 Y vdd vss
** Your code **
.ends

…